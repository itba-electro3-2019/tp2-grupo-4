module Gen_Com(out);
    output out;
    assign out=1;
endmodule