module In(out);
    output [4:0] out;
    assign out=5'b01001;
endmodule